module UART_Tx();





endmodule 
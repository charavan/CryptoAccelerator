module Testbench;




endmodule 
module UART_Rx();




endmodule 
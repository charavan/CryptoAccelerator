module Maj( input  [31:0] a , b , c ,
            output [31:0]            out1,out2);




assign out = (a & b) | (c & (a | b) );

endmodule 
module T_two ( input  [31:0] s0, maj ,
               output [31:0] out      );



assign out = s0 + maj ;



endmodule 